module tb_ula_74181;

logic[3:0] a, b, s;
logic m, c_in;

ula_74181 uut(.a());

initial
begin
    
    
    $stop;
end
endmodule